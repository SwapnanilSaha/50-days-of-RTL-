module clock(clk_in);
input clk_in;
endmodule

