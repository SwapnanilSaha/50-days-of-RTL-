module receiver_tb;
reg [47:0]d;
wire out;
receiver v1(d,out);
initial
begin
d= 48'b100111010010110111000011110101011001111011111100;
#5;
d= 48'b100111010010110111000011110101011001111011111101;
#5;
d=48'b100111010010110111100111110101011001111011111100;
#5;
 d=48'b100111010010110111000011110101011001111011111100;
#5 $finish;
end
endmodule
